library verilog;
use verilog.vl_types.all;
entity multiplexador_vlg_vec_tst is
end multiplexador_vlg_vec_tst;
