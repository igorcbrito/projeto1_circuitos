library verilog;
use verilog.vl_types.all;
entity tratamentoSubtracao_vlg_vec_tst is
end tratamentoSubtracao_vlg_vec_tst;
