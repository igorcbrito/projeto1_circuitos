library verilog;
use verilog.vl_types.all;
entity menorque_vlg_vec_tst is
end menorque_vlg_vec_tst;
